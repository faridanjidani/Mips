module ALU(
	input [31:0] in1,
	input [31:0] in2,
	input [3:0] cmd,
	output reg [31:0] result
	);

	always @(*) begin
		case (cmd)
			4'b0000: result = in1 + in2;

			4'b0010: result = in1 - in2;

			4'b0100: result = in1 & in2;

			4'b0101: result = in1 | in2;

			4'b0110: result = ~ (in1 | in2);

			4'b0111: result = in1 ^ in2;

			4'b1000: result = in1 << in2;

			4'b1001:
			begin
				// result = in1 >>> in2;  // system verilog
	      		case(in2)
	      			0:  result = in1;
	      			1:  result = in1[31] == 1'b1 ? {1'b1, in1[31:1]}  : {1'b0, in1[31:1]};
	      			2:  result = in1[31] == 1'b1 ? {2'b11, in1[31:2]}  : {2'b0, in1[31:2]};
	      			3:  result = in1[31] == 1'b1 ? {3'b111, in1[31:3]}  : {3'b0, in1[31:3]};
	      			4:  result = in1[31] == 1'b1 ? {4'b1111, in1[31:4]}  : {4'b0, in1[31:4]};
	      			5:  result = in1[31] == 1'b1 ? {5'b11111, in1[31:5]}  : {5'b0, in1[31:5]};
	      			6:  result = in1[31] == 1'b1 ? {6'b111111, in1[31:6]}  : {6'b0, in1[31:6]};
	      			7:  result = in1[31] == 1'b1 ? {7'b1111111, in1[31:7]}  : {7'b0, in1[31:7]};
	      			8:  result = in1[31] == 1'b1 ? {8'b11111111, in1[31:8]}  : {8'b0, in1[31:8]};
	      			9:  result = in1[31] == 1'b1 ? {9'b111111111, in1[31:9]}  : {9'b0, in1[31:9]};
	      			10: result = in1[31] == 1'b1 ? {10'b1111111111, in1[31:10]} : {10'b0, in1[31:10]};
	      			11: result = in1[31] == 1'b1 ? {11'b11111111111, in1[31:11]} : {11'b0, in1[31:11]};
	      			12: result = in1[31] == 1'b1 ? {12'b111111111111, in1[31:12]} : {12'b0, in1[31:12]};
	      			13: result = in1[31] == 1'b1 ? {13'b1111111111111, in1[31:13]} : {13'b0, in1[31:13]};
	      			14: result = in1[31] == 1'b1 ? {14'b11111111111111, in1[31:14]} : {14'b0, in1[31:14]};
	      			15: result = in1[31] == 1'b1 ? {15'b111111111111111, in1[31:15]} : {15'b0, in1[31:15]};
	      			16: result = in1[31] == 1'b1 ? {16'b1111111111111111, in1[31:16]} : {16'b0, in1[31:16]};
	      			17: result = in1[31] == 1'b1 ? {17'b11111111111111111, in1[31:17]} : {17'b0, in1[31:17]};
	      			18: result = in1[31] == 1'b1 ? {18'b111111111111111111, in1[31:18]} : {18'b0, in1[31:18]};
	      			19: result = in1[31] == 1'b1 ? {19'b1111111111111111111, in1[31:19]} : {19'b0, in1[31:19]};
	      			20: result = in1[31] == 1'b1 ? {20'b11111111111111111111, in1[31:20]} : {20'b0, in1[31:20]};
	      			21: result = in1[31] == 1'b1 ? {21'b111111111111111111111, in1[31:21]} : {21'b0, in1[31:21]};
	      			22: result = in1[31] == 1'b1 ? {22'b1111111111111111111111, in1[31:22]}  : {22'b0, in1[31:22]};
	      			23: result = in1[31] == 1'b1 ? {23'b11111111111111111111111, in1[31:23]}  : {23'b0, in1[31:23]};
	      			24: result = in1[31] == 1'b1 ? {24'b111111111111111111111111, in1[31:24]}  : {24'b0, in1[31:24]};
	      			25: result = in1[31] == 1'b1 ? {25'b1111111111111111111111111, in1[31:25]}  : {25'b0, in1[31:25]};
	      			26: result = in1[31] == 1'b1 ? {26'b11111111111111111111111111, in1[31:26]}  : {26'b0, in1[31:26]};
	      			27: result = in1[31] == 1'b1 ? {27'b111111111111111111111111111, in1[31:27]}  : {27'b0, in1[31:27]};
	      			28: result = in1[31] == 1'b1 ? {28'b1111111111111111111111111111, in1[31:28]}  : {28'b0, in1[31:28]};
	      			29: result = in1[31] == 1'b1 ? {29'b11111111111111111111111111111, in1[31:29]}  : {29'b0, in1[31:29]};
	      			30: result = in1[31] == 1'b1 ? {30'b111111111111111111111111111111, in1[31:30]}  : {30'b0, in1[31:30]};
	      			31: result = in1[31] == 1'b1 ? {31'b1111111111111111111111111111111, in1[31]}    : {31'b0, in1[31]};
	      		endcase
	      	end
			4'b1010: result = in1 >> in2;

			default: result = in1 + in2;
		endcase
	end

endmodule